module tt_slave (
input 			req,
input [31:0]	addr,
input 			cmd,
input [31:0]	wdata,
output 			ack,
output [31:0]	rdata
);










endmodule