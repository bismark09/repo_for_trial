module tt_tb();


tt_crossbar #(2,2)(

input 			master_req 		[NUM_MASTER-1],
input [31:0]	master_addr 	[NUM_MASTER-1],
input 			master_cmd		[NUM_MASTER-1],
input [31:0]	master_wdata	[NUM_MASTER-1],
output 			master_ack		[NUM_MASTER-1],
output [31:0]	master_rdata	[NUM_MASTER-1],


);






endmodule