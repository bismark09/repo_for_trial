module cross_bar(



);



endmodule 