
interface tt_bus_irf(
	logic 			req,
	logic [31:0]	addr,
	logic 			cmd,
	logic [31:0]	wdata,
	logic 			ack,
	logic [31:0]	rdata
);


endinterface
