module tt_tb();




endmodule