module tt_crossbar(



);



endmodule 