module tt_slave (
output 			req,
output [31:0]	addr,
output 			cmd,
output [31:0]	wdata,
input 			ack,
input  [31:0]	rdata
);



endmodule